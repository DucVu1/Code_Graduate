library verilog;
use verilog.vl_types.all;
entity matching_stage_vlg_vec_tst is
end matching_stage_vlg_vec_tst;
